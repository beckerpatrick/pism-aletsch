netcdf pism_overrides {
    variables:
    byte pism_overrides;

   pism_overrides:run_title = "PISM Aletschgletscher";
   pism_overrides:run_title_doc = "Free-form string containing a concise description of the current run. This string is written to output files as the 'title' global attribute.";

    pism_overrides:bed_smoother_range = 0.;
    pism_overrides:bed_smoother_range_doc = "m; half-width of smoothing domain for PISMBedSmoother, in implementing [\\ref Schoofbasaltopg2003] bed roughness parameterization for SIA; set value to zero to turn off mechanism";

    pism_overrides:summary_vol_scale_factor_log10 = 0;
    pism_overrides:summary_vol_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for volume (in km^3) in summary line to stdout";

    pism_overrides:summary_area_scale_factor_log10 = 0;
    pism_overrides:summary_area_scale_factor_log10_doc = "; an integer; log base 10 of scale factor to use for area (in km^2) in summary line to stdout";

    pism_overrides:ice_softness = 2.25e-24;
    pism_overrides:ice_softness_doc = "Pa-3 s-1; ice softness used by IsothermalGlenIce";

    pism_overrides:pseudo_plastic_uthreshold = 50.0;
    pism_overrides:pseudo_plastic_uthreshold_doc = "m/year; ";

}